module new( 
    input x, 
    output y
);

    always @(x) begin end

    assign y = 1;
endmodule