`ifndef __TIMESCALE_VH__
`define __TIMESCALE_VH__

`timescale 1ns/1ps

`endif // __TIMESCALE_VH__