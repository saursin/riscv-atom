///////////////////////////////////////////////////////////////////
//  File        : Timescale.vh
//  Author      : Saurabh Singh (saurabh.s99100@gmail.com)
//  Description : Timescale header file
///////////////////////////////////////////////////////////////////

`ifndef __TIMESCALE_VH__
`define __TIMESCALE_VH__

`timescale 1ns/1ps

`endif // __TIMESCALE_VH__
