`default_nettype none

module spi
(
    
);

endmodule